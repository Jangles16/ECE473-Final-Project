//IF_ID_pipe.v

module IF_ID_pipe(
	input wire clock,
	input wire [31:0] PC_in,
	input wire [31:0] instr_in,
	output reg [31:0] PC_out,
	output reg [31:0]	instr_out
	);
	
	
	always @(posedge clock) begin
		PC_out<=PC_in;
		instr_out<=instr_in;
	end
endmodule