//char_engine
//version 2 (in progress)
//changed from previous: extending the character set to support the full alphabet, and special characters

//This character display enginne is designed to work with CPU developement projects, and displays various information from the project onto a vga-monitor.
//There is a built in hex engine that runs off the 3 data sources from the project.
//Characters are 8 * 8 pixels each with a blank line above each character, allowing allowing 80 * 53 characters on screen.
//The memory mapping takes into account only a 640*480 screen resolution

module char_engine(
	input wire clock,
	input wire project_clock,

	input wire [31:0] ins_data, //these inputs are for the data to be displayed later
	input wire [31:0] mem_data,
	input wire [31:0] reg_data,
	input wire [15:0] prg_counter,
	input wire [15:0]	cycle_counter,
	input wire [31:0] debug, //debug input
	input wire [31:0] gp_reg_1, //General Purpose Register inputs
	input wire [31:0] gp_reg_2,
	input wire [31:0] gp_reg_3,
	input wire [31:0] gp_reg_4,
	input wire [31:0] gp_reg_5, //General Purpose Register inputs
	input wire [31:0] gp_reg_6,
	input wire [31:0] gp_reg_7,
	input wire [31:0] gp_reg_8,	
	
	output reg [0:7] mem_out, //if everything is backwards, swap the bit order on this output and recompile!
	output reg [15:0] mem_add,
	output mem_write,
	
	output reg [4:0] reg_sw,
	output reg [5:0] ins_sw,
	output reg [5:0] mem_sw);
	
	assign mem_write = 1;
	
	reg [6:0] hex_digit;
	reg [31:0] data;
	reg [5:0] hex_buffer[0:(MAX_STRING_LENGTH - 1)];
	reg [5:0] debug_prebuffer[0:31];
	reg [5:0] debug_buffer[0:38];
	reg [15:0] pc_history[0:9];
	reg [63:0] mem_buffer;
	
	parameter HORI_OFFSET = 0; //sets the horizontal offset of the memory renderer, only use if the top of the screen gets cut off.
	parameter NUM_LABEL_TASKS = 20; // This tells the code where to start tasks that require data manipulation, this must be set as you add more labels, debug tasks must be part of this number
	parameter MAX_STRING_LENGTH = 20; //Generally you do not need to modify this, but it will change the global maximum string length (default = 20)
	parameter DEBUG_TRUE = 6'h01; //This will change the charcter used when a debug value comes back as true
	parameter DEBUG_FALSE = 6'h00; //This will change the character used when a debug value comes back as false
	
	
	
	integer debug_count;
	
	integer data_index, reg_index, row, column, slice_delay, decode_delay, num_chars, k, x, y, z;
	
	initial begin
	slice_delay = 0; //initial values for the character renderer
	decode_delay = 0;
	x = 0;
	y = -1;
	data_index = -1;
	reg_index = 0;
	debug_count = 0;
	end
	
	always @(posedge clock) begin //semi-pipelined design, only executes one if statement per clock
				
		if (x < 0) begin //source and slice steps
			if (slice_delay == 0) data_index = data_index + 1;
			source_data();
			if (data_index > NUM_LABEL_TASKS) slice_data ();
			slice_delay = slice_delay + 1;
			if (slice_delay == 2) begin
				x = num_chars - 1;
				slice_delay = 0;
			end
		end
		
		else if (y < 0) begin //decode steps
			hex_digit <= hex_buffer[x];
			if (decode_delay == 0) begin
				x = x - 1;
			end
			decode_hex();
			decode_delay = decode_delay + 1;
			if (decode_delay == 3) begin
				y = 8;
				decode_delay = 0;
			end
		end
		
		else if (y >= 0) begin //this step writes to memory
			k = (y * 8) - 1;
			mem_add <= (80 * y) + (800 * row) + (num_chars - (x + 1)) + (column) + (HORI_OFFSET * 80); //this complicated formula tranlates information into a linear address
			mem_out <= mem_buffer[k -: 8];
			y = y - 1;
		end
	end
	
	always @(posedge clock) begin //debug indicators are set here
		
		if (debug[debug_count] == 1) debug_prebuffer[debug_count] <= DEBUG_TRUE; //this is the printed character for a true result, default = T
		else debug_prebuffer[debug_count] <= DEBUG_FALSE; //this is the character printed for a false result, default = F
		debug_count = debug_count + 1;
		if (debug_count > 31) debug_count = 0;
	end
	
	always @(posedge project_clock) begin //the program counter history is set by this code, it is driven by the clock of the project so that the data does not update too fast
		if (prg_counter != pc_history[0]) begin
			pc_history[9] = pc_history[8];
			pc_history[8] = pc_history[7];
			pc_history[7] = pc_history[6];
			pc_history[6] = pc_history[5];
			pc_history[5] = pc_history[4];
			pc_history[4] = pc_history[3];
			pc_history[3] = pc_history[2];
			pc_history[2] = pc_history[1];
			pc_history[1] = pc_history[0];
			pc_history[0] = prg_counter;
		end
	end
	always begin 
	//this is brute force way of building the debug buffer with spaces in it, the other methods used more logic units, and did not work properly due to timing issues
	//this method uses constant assignment to build the proper string, which uses far fewer LUs.	
	// I tried doing this procedurely using a loop, but found that it ran into timing issues, so I just use the direct method.
		debug_buffer[0] = 6'h24;
		debug_buffer[1] = debug_prebuffer[0];
		debug_buffer[2] = debug_prebuffer[1];
		debug_buffer[3] = debug_prebuffer[2];
		debug_buffer[4] = debug_prebuffer[3];
		debug_buffer[5] = 6'h24;
		debug_buffer[6] = debug_prebuffer[4];
		debug_buffer[7] = debug_prebuffer[5];
		debug_buffer[8] = debug_prebuffer[6];
		debug_buffer[9] = debug_prebuffer[7];
		debug_buffer[10] = 6'h24;
		debug_buffer[11] = debug_prebuffer[8];
		debug_buffer[12] = debug_prebuffer[9];
		debug_buffer[13] = debug_prebuffer[10];
		debug_buffer[14] = debug_prebuffer[11];
		debug_buffer[15] = 6'h24;
		debug_buffer[16] = debug_prebuffer[12];
		debug_buffer[17] = debug_prebuffer[13];
		debug_buffer[18] = debug_prebuffer[14];
		debug_buffer[19] = debug_prebuffer[15];
		debug_buffer[20] = debug_prebuffer[16];
		debug_buffer[21] = debug_prebuffer[17];
		debug_buffer[22] = debug_prebuffer[18];
		debug_buffer[23] = debug_prebuffer[19];
		debug_buffer[24] = 6'h24;
		debug_buffer[25] = debug_prebuffer[20];
		debug_buffer[26] = debug_prebuffer[21];
		debug_buffer[27] = debug_prebuffer[22];
		debug_buffer[28] = debug_prebuffer[23];
		debug_buffer[29] = 6'h24;
		debug_buffer[30] = debug_prebuffer[24];
		debug_buffer[31] = debug_prebuffer[25];
		debug_buffer[32] = debug_prebuffer[26];
		debug_buffer[33] = debug_prebuffer[27];
		debug_buffer[34] = 6'h24;
		debug_buffer[35] = debug_prebuffer[28];
		debug_buffer[36] = debug_prebuffer[29];
		debug_buffer[37] = debug_prebuffer[30];
		debug_buffer[38] = debug_prebuffer[31];
	end
	
	task source_data; //This part of the module is the main task list for the renderer, it can be utilized in a variety of ways to render information.
			
		if (data_index == NUM_LABEL_TASKS + 4) ins_sw <= reg_index;
		if (data_index == NUM_LABEL_TASKS + 5) ins_sw <= reg_index + 32; //this code requests the data from memory to be printed on screen
		if (data_index == NUM_LABEL_TASKS + 6) mem_sw <= reg_index;
		if (data_index == NUM_LABEL_TASKS + 7) mem_sw <= reg_index + 32; //it always request the data one clock ahead of time, so that the data is ready when the system reads it
		// Two lines below added by Nicholas LaJoie - corrects register data formatting on screen
		if (data_index == NUM_LABEL_TASKS + 8) reg_sw <= reg_index; 
		//if (data_index == NUM_LABEL_TASKS + 9) reg_sw <= reg_index + 32; //this line is not needed, as there are only 32 registers
		
		case (data_index)
		//in the case of text labels, the hex_buffer is set manually for each character, and the data is only written to memory once.
			0: begin //"INS. MEMORY" label
				hex_buffer[10] <= 6'h12;
				hex_buffer[9] <= 6'h17;
				hex_buffer[8] <= 6'h1C;
				hex_buffer[7] <= 6'h28;
				hex_buffer[6] <= 6'h24;
				hex_buffer[5] <= 6'h16;
				hex_buffer[4] <= 6'h0E;
				hex_buffer[3] <= 6'h16;
				hex_buffer[2] <= 6'h18;
				hex_buffer[1] <= 6'h1B;
				hex_buffer[0] <= 6'h22;
				
				row = 0;
				column = 0;
				num_chars = 11;
				end
			
			1: begin //"DATA MEMORY" label
					hex_buffer[10] <= 6'h0D;
					hex_buffer[9] <= 6'h0A;
					hex_buffer[8] <= 6'h1D;
					hex_buffer[7] <= 6'h0A;
					hex_buffer[6] <= 6'h24;
					hex_buffer[5] <= 6'h16;
					hex_buffer[4] <= 6'h0E;
					hex_buffer[3] <= 6'h16;
					hex_buffer[2] <= 6'h18;
					hex_buffer[1] <= 6'h1B;
					hex_buffer[0] <= 6'h22;
					
					row = 0;
					column = 25;
					num_chars = 11;
				end
				
			2: begin //"REGISTERS" label
					hex_buffer[8] <= 6'h1B;
					hex_buffer[7] <= 6'h0E;
					hex_buffer[6] <= 6'h10;
					hex_buffer[5] <= 6'h12;
					hex_buffer[4] <= 6'h1C;
					hex_buffer[3] <= 6'h1D;
					hex_buffer[2] <= 6'h0E;
					hex_buffer[1] <= 6'h1B;
					hex_buffer[0] <= 6'h1C;
					
					row = 0;
					column = 50;
					num_chars = 9;
				end
				
				3: begin //PC HISTORY label
						hex_buffer[9] <= 6'h19;
						hex_buffer[8] <= 6'h0C;
						hex_buffer[7] <= 6'h24;
						hex_buffer[6] <= 6'h11;
						hex_buffer[5] <= 6'h12;
						hex_buffer[4] <= 6'h1C;
						hex_buffer[3] <= 6'h1D;
						hex_buffer[2] <= 6'h18;
						hex_buffer[1] <= 6'h1B;
						hex_buffer[0] <= 6'h22;			
					
						row  = 0;
						column = 63;
						num_chars = 10;
					end
					
				4: begin //CYCLES label
						hex_buffer[6] <= 6'h0C;
						hex_buffer[5] <= 6'h22;
						hex_buffer[4] <= 6'h0C;
						hex_buffer[3] <= 6'h15;
						hex_buffer[2] <= 6'h0E;
						hex_buffer[1] <= 6'h1C;
						hex_buffer[0] <= 6'h27;
				
						row = 35;
						column = 0;
						num_chars = 7;
					end
				5: begin //DEBUG label
						hex_buffer[4] <= 6'h0D;
						hex_buffer[3] <= 6'h0E;
						hex_buffer[2] <= 6'h0B;
						hex_buffer[1] <= 6'h1E;
						hex_buffer[0] <= 6'h10;
				
						row = 39;
						column = 0;
						num_chars = 5;
					end
					
				6: begin //Current PC
						
						hex_buffer[9] <= 6'h0c;
						hex_buffer[8] <= 6'h1e;
						hex_buffer[7] <= 6'h1b;
						hex_buffer[6] <= 6'h1b;
						hex_buffer[5] <= 6'h0e;
						hex_buffer[4] <= 6'h17;
						hex_buffer[3] <= 6'h1d;
						hex_buffer[2] <= 6'h24;
						hex_buffer[1] <= 6'h19;
						hex_buffer[0] <= 6'h0c;
						
						row = 13;
						column = 63;
						num_chars = 10;
					end
					
				7: begin //IF ID INSTR
						
						hex_buffer[10] <= 6'h12;
						hex_buffer[9] <= 6'h0f;
						hex_buffer[8] <= 6'h24;
						hex_buffer[7] <= 6'h12;
						hex_buffer[6] <= 6'h0d;
						hex_buffer[5] <= 6'h24;
						hex_buffer[4] <= 6'h12;
						hex_buffer[3] <= 6'h17;
						hex_buffer[2] <= 6'h1c;
						hex_buffer[1] <= 6'h1d;
						hex_buffer[0] <= 6'h1b;
						
						row = 16;
						column = 63;
						num_chars = 11;
					end
					
				8: begin //Branch Addr
						
						hex_buffer[10] <= 6'h0b;
						hex_buffer[9] <= 6'h1b;
						hex_buffer[8] <= 6'h0a;
						hex_buffer[7] <= 6'h17;
						hex_buffer[6] <= 6'h0c;
						hex_buffer[5] <= 6'h11;
						hex_buffer[4] <= 6'h24;
						hex_buffer[3] <= 6'h0a;
						hex_buffer[2] <= 6'h0d;
						hex_buffer[1] <= 6'h0d;
						hex_buffer[0] <= 6'h1b;
						
						row = 19;
						column = 63;
						num_chars = 11;
					end
			
				9: begin //EX MEM FW
					
						hex_buffer[8] <= 6'h0e;
						hex_buffer[7] <= 6'h21;
						hex_buffer[6] <= 6'h24;
						hex_buffer[5] <= 6'h16;
						hex_buffer[4] <= 6'h0e;
						hex_buffer[3] <= 6'h16;
						hex_buffer[2] <= 6'h24;
						hex_buffer[1] <= 6'h0f;
						hex_buffer[0] <= 6'h20;
						
						row = 22;
						column = 63;
						num_chars = 9;
					end
					

				10: begin //RAM OUT
						
						hex_buffer[6] <= 6'h1b;
						hex_buffer[5] <= 6'h0a;
						hex_buffer[4] <= 6'h16;
						hex_buffer[3] <= 6'h24;
						hex_buffer[2] <= 6'h18;
						hex_buffer[1] <= 6'h1e;
						hex_buffer[0] <= 6'h1d;
						
						row = 25;
						column = 63;
						num_chars = 7;
					end

				11: begin //RAM WRITE
						
						hex_buffer[8] <= 6'h1b;
						hex_buffer[7] <= 6'h0a;
						hex_buffer[6] <= 6'h16;
						hex_buffer[5] <= 6'h24;
						hex_buffer[4] <= 6'h20;
						hex_buffer[3] <= 6'h1b;
						hex_buffer[2] <= 6'h12;
						hex_buffer[1] <= 6'h1d;
						hex_buffer[0] <= 6'h0e;
						
						row = 28;
						column = 63;
						num_chars = 9;
					end

				12: begin //WRITE DATA
						
						hex_buffer[9] <= 6'h20;
						hex_buffer[8] <= 6'h1b;
						hex_buffer[7] <= 6'h12;
						hex_buffer[6] <= 6'h1d;
						hex_buffer[5] <= 6'h0e;
						hex_buffer[4] <= 6'h24;
						hex_buffer[3] <= 6'h0d;
						hex_buffer[2] <= 6'h0a;
						hex_buffer[1] <= 6'h1d;
						hex_buffer[0] <= 6'h0a;
						
						row = 31;
						column = 63;
						num_chars = 10;
					end

				13: begin //WRITE ADDR
						
						hex_buffer[9] <= 6'h20;
						hex_buffer[8] <= 6'h1b;
						hex_buffer[7] <= 6'h12;
						hex_buffer[6] <= 6'h1d;
						hex_buffer[5] <= 6'h0e;
						hex_buffer[4] <= 6'h24;
						hex_buffer[3] <= 6'h0a;
						hex_buffer[2] <= 6'h0d;
						hex_buffer[1] <= 6'h0d;
						hex_buffer[0] <= 6'h1b;
						
						row = 34;
						column = 63;
						num_chars = 10;
					end					
					
				14: begin //00-15: label
						hex_buffer[5] <= 6'h00;
						hex_buffer[4] <= 6'h00;
						hex_buffer[3] <= 6'h26;
						hex_buffer[2] <= 6'h01;
						hex_buffer[1] <= 6'h05;
						hex_buffer[0] <= 6'h27;
						
						row = 40;
						column = 0;
						num_chars = 6;
					end
				15: begin //16-31: label
						hex_buffer[5] <= 6'h01;
						hex_buffer[4] <= 6'h06;
						hex_buffer[3] <= 6'h26;
						hex_buffer[2] <= 6'h03;
						hex_buffer[1] <= 6'h01;
						hex_buffer[0] <= 6'h27;
					
						row = 42;
						column = 0;
						num_chars = 6;
					end
				
				16: begin //debug 0-15 task
					z = 0;
				
					while (z <= 19) begin
						hex_buffer[z] = debug_buffer[z];
						z = z + 1;
					end
					
					column = 6;
					row = 40;
					num_chars = 20;
				end
				
			17: begin //debug 16-31 task
					z = 0;
				
					while (z <= 18) begin
						hex_buffer[z] = debug_buffer[z + 20];
						z = z + 1;
					end
					
					column = 6;
					row = 42;
					num_chars = 19;
				end
				
				
/******************************************************

******************CHANGE THIS STUFF********************

*******************************************************/	

			
			18: begin //just my name
			
					hex_buffer[11] <= 6'h13;
					hex_buffer[10] <= 6'h18;
					hex_buffer[9] <= 6'h1c;
					hex_buffer[8] <= 6'h11;
					hex_buffer[7] <= 6'h24;
					hex_buffer[6] <= 6'h0a;
					hex_buffer[5] <= 6'h17;
					hex_buffer[4] <= 6'h0d;
					hex_buffer[3] <= 6'h1b;
					hex_buffer[2] <= 6'h0e;
					hex_buffer[1] <= 6'h20;
					hex_buffer[0] <= 6'h1c;
					
					row = 40;
					column = 50;
					num_chars = 12;
			end
			
			19: begin //milestone #
			
					hex_buffer[10] <= 6'h16;
					hex_buffer[9] <= 6'h12;
					hex_buffer[8] <= 6'h15;
					hex_buffer[7] <= 6'h0e;
					hex_buffer[6] <= 6'h1c;
					hex_buffer[5] <= 6'h1d;
					hex_buffer[4] <= 6'h18;
					hex_buffer[3] <= 6'h17;
					hex_buffer[2] <= 6'h0e;
					hex_buffer[1] <= 6'h24;
					hex_buffer[0] <= 6'h04;		//change to hex # of current milestone
					
					row = 41;
					column = 50;
					num_chars = 11;
			end
			
			20: begin // Test #
			
					hex_buffer[5] <= 6'h1d;
					hex_buffer[4] <= 6'h0e;
					hex_buffer[3] <= 6'h1c;
					hex_buffer[2] <= 6'h1d;
					hex_buffer[1] <= 6'h24;
					hex_buffer[0] <= 6'h05;		//change to hex number of current test
					
					row = 42;
					column = 50;
					num_chars = 6;
			end
			(NUM_LABEL_TASKS + 1): begin //instruction memory indexes 00-31
					data <= reg_index;
					column = 0;
					row = reg_index + 1;
					num_chars = 2;
				end
			
			(NUM_LABEL_TASKS + 2): begin //instruction memory indexes 32-63
					data <= reg_index + 32;
					column = 12;
					row = reg_index + 1;
					num_chars = 2;
				end	
				
			(NUM_LABEL_TASKS + 3): begin //data_memory indexes 00-31
					data <= reg_index;
					column = 25;
					row = reg_index + 1;
					num_chars = 2;
				end
				
			(NUM_LABEL_TASKS + 4): begin //data_memory indexes 32-63
					data <= reg_index + 32;
					column = 37;
					row = reg_index + 1;
					num_chars = 2;
				end
				
			(NUM_LABEL_TASKS + 5): begin //instruction memory data 00-31
					data <= ins_data;
					column = 2;
					row = reg_index + 1;
					num_chars = 9;
					hex_buffer[8] <= 6'h27;
				end
				
			(NUM_LABEL_TASKS + 6): begin //instruction memory data 32-63
					data <= ins_data;
					column = 14;
					row = reg_index + 1;
					num_chars = 9;
					hex_buffer[8] <= 6'h27;
				end
			
			(NUM_LABEL_TASKS + 7): begin //data memory data 00-31
					data <= mem_data; 
					column = 27;
					row = reg_index + 1;
					num_chars = 9;
					hex_buffer[8] <= 6'h27;
				end
			
			(NUM_LABEL_TASKS + 8): begin //data memory data 31-63
					data <= mem_data; 
					column = 39;
					row = reg_index + 1;
					num_chars = 9;
					hex_buffer[8] <= 6'h27;
				end
				
			(NUM_LABEL_TASKS + 9): begin //register indexes
					data <= 0;
					data[4:0] <= reg_index;
					column = 50;
					row = reg_index + 1;
					num_chars = 2;
				end
				
			(NUM_LABEL_TASKS + 10): begin // register data
					reg_sw <= reg_index;
					data <= reg_data;
					column = 52;
					row = reg_index + 1;
					num_chars = 9;
					hex_buffer[8] <= 6'h27;
					if (slice_delay == 1) reg_index = reg_index + 1;
					if (reg_index == 32) begin //this resets the register index variable to zero once it reaches 32
						reg_index = 0;
					end
				end
			
			(NUM_LABEL_TASKS + 11): begin //Cycles data
					data <= cycle_counter; 
					column = 8;
					row = 35;
					num_chars = 4;
				end
			
			(NUM_LABEL_TASKS + 12): begin //pc history data
					if (reg_index <= 9) begin
						data <= pc_history[reg_index];
						row = reg_index + 1;
						column = 63;
						num_chars = 4;
					end
				
					else num_chars = 0; //setting num chars to 0 causes nothing to be written to memory, essentially aborting the source_data task
				
				end 
			(NUM_LABEL_TASKS + 13): begin
					data <= gp_reg_1;
					column = 63;
					row = 14;
					num_chars = 8;
				end
		
			(NUM_LABEL_TASKS + 14): begin
					data <= gp_reg_2;
					column = 63;
					row = 17;
					num_chars = 8;
				end
				
			(NUM_LABEL_TASKS + 15): begin
					data <= gp_reg_3;
					column = 63;
					row = 20;
					num_chars = 8;
				end

			(NUM_LABEL_TASKS + 16): begin
					data <= gp_reg_4;
					column = 63;
					row = 23;
					num_chars = 8;
				end
				

			(NUM_LABEL_TASKS + 17): begin
					data <= gp_reg_5;
					column = 63;
					row = 26;
					num_chars = 8;
				end

			(NUM_LABEL_TASKS + 18): begin
					data <= gp_reg_6;
					column = 63;
					row = 29;
					num_chars = 8;
				end

			(NUM_LABEL_TASKS + 19): begin
					data <= gp_reg_7;
					column = 63;
					row = 32;
					num_chars = 8;
				end

			(NUM_LABEL_TASKS + 20): begin
					data <= gp_reg_8;
					column = 63;
					row = 35;
					num_chars = 8;
				end
				
			default: data_index = NUM_LABEL_TASKS;
		endcase
	endtask
	
	task slice_data; //I tried other ways of doing this, but the straightforward approach works better.
		hex_buffer[7] <= data[31:28];
		hex_buffer[6] <= data[27:24];
		hex_buffer[5] <= data[23:20];
		hex_buffer[4] <= data[19:16];
		hex_buffer[3] <= data[15:12];
		hex_buffer[2] <= data[11:8];
		hex_buffer[1] <= data[7:4];
		hex_buffer[0] <= data[3:0];
	endtask
	
	task decode_hex;
		case (hex_digit)	
		
			6'h00: begin //zero
					mem_buffer[7:0] <=   8'b00111100;
					mem_buffer[15:8] <=  8'b01000010;
					mem_buffer[23:16] <= 8'b01000010;
					mem_buffer[31:24] <= 8'b01000010;
					mem_buffer[39:32] <= 8'b01000010;
					mem_buffer[47:40] <= 8'b01000010;
					mem_buffer[55:48] <= 8'b01000010;
					mem_buffer[63:56] <= 8'b00111100;
					end
			
			6'h01: begin //one
					mem_buffer[7:0] <=   8'b00011000;
					mem_buffer[15:8] <=  8'b00111000;
					mem_buffer[23:16] <= 8'b01111000;
					mem_buffer[31:24] <= 8'b00011000;
					mem_buffer[39:32] <= 8'b00011000;
					mem_buffer[47:40] <= 8'b00011000;
					mem_buffer[55:48] <= 8'b00011000;
					mem_buffer[63:56] <= 8'b01111110;
					end
			
			6'h02: begin //two
					mem_buffer[7:0] <=   8'b00111100;
					mem_buffer[15:8] <=  8'b01100110;
					mem_buffer[23:16] <= 8'b01100110;
					mem_buffer[31:24] <= 8'b00001100;
					mem_buffer[39:32] <= 8'b00011000;
					mem_buffer[47:40] <= 8'b00110000;
					mem_buffer[55:48] <= 8'b01100000;
					mem_buffer[63:56] <= 8'b01111110;
					end
					
			6'h03: begin //three
					mem_buffer[7:0] <=   8'b01111100;
					mem_buffer[15:8] <=  8'b00000110;
					mem_buffer[23:16] <= 8'b00000110;
					mem_buffer[31:24] <= 8'b01111100;
					mem_buffer[39:32] <= 8'b00000110;
					mem_buffer[47:40] <= 8'b00000110;
					mem_buffer[55:48] <= 8'b00000110;
					mem_buffer[63:56] <= 8'b01111100;
					end
				
			6'h04: begin //four
					mem_buffer[7:0] <=   8'b00001110;
					mem_buffer[15:8] <=  8'b00010110;
					mem_buffer[23:16] <= 8'b00100110;
					mem_buffer[31:24] <= 8'b01000110;
					mem_buffer[39:32] <= 8'b01000110;
					mem_buffer[47:40] <= 8'b01111110;
					mem_buffer[55:48] <= 8'b00000110;
					mem_buffer[63:56] <= 8'b00000110;
					end
					
			6'h05: begin //five
					mem_buffer[7:0] <=   8'b01111110;
					mem_buffer[15:8] <=  8'b01100000;
					mem_buffer[23:16] <= 8'b01100000;
					mem_buffer[31:24] <= 8'b01111000;
					mem_buffer[39:32] <= 8'b00001100;
					mem_buffer[47:40] <= 8'b00000110;
					mem_buffer[55:48] <= 8'b00001100;
					mem_buffer[63:56] <= 8'b01111000;
					end
					
			6'h06: begin //six
					mem_buffer[7:0] <=   8'b00111100;
					mem_buffer[15:8] <=  8'b01000000;
					mem_buffer[23:16] <= 8'b01000000;
					mem_buffer[31:24] <= 8'b01111100;
					mem_buffer[39:32] <= 8'b01000010;
					mem_buffer[47:40] <= 8'b01000010;
					mem_buffer[55:48] <= 8'b01000010;
					mem_buffer[63:56] <= 8'b00111100;
					end
					
			6'h07: begin //seven
					mem_buffer[7:0] <=   8'b01111110;
					mem_buffer[15:8] <=  8'b00000110;
					mem_buffer[23:16] <= 8'b00000110;
					mem_buffer[31:24] <= 8'b00000110;
					mem_buffer[39:32] <= 8'b00001100;
					mem_buffer[47:40] <= 8'b00011000;
					mem_buffer[55:48] <= 8'b00110000;
					mem_buffer[63:56] <= 8'b01100000;
					end
					
			6'h08: begin //eight
					mem_buffer[7:0] <=   8'b00111100;
					mem_buffer[15:8] <=  8'b01000010;
					mem_buffer[23:16] <= 8'b01000010;
					mem_buffer[31:24] <= 8'b00111100;
					mem_buffer[39:32] <= 8'b01000010;
					mem_buffer[47:40] <= 8'b01000010;
					mem_buffer[55:48] <= 8'b01000010;
					mem_buffer[63:56] <= 8'b00111100;
					end
					
			6'h09: begin //nine
					mem_buffer[7:0] <=   8'b00111100;
					mem_buffer[15:8] <=  8'b01000110;
					mem_buffer[23:16] <= 8'b01000110;
					mem_buffer[31:24] <= 8'b01000110;
					mem_buffer[39:32] <= 8'b00111110;
					mem_buffer[47:40] <= 8'b00000110;
					mem_buffer[55:48] <= 8'b00000110;
					mem_buffer[63:56] <= 8'b00000110;
					end
					
			6'h0A: begin //A
					mem_buffer[7:0] <=   8'b00111100;
					mem_buffer[15:8] <=  8'b01000010;
					mem_buffer[23:16] <= 8'b01000010;
					mem_buffer[31:24] <= 8'b01000010;
					mem_buffer[39:32] <= 8'b01111110;
					mem_buffer[47:40] <= 8'b01000010;
					mem_buffer[55:48] <= 8'b01000010;
					mem_buffer[63:56] <= 8'b01000010;
					end
					
			6'h0B: begin //B
					mem_buffer[7:0] <=   8'b01111100;
					mem_buffer[15:8] <=  8'b01000010;
					mem_buffer[23:16] <= 8'b01000110;
					mem_buffer[31:24] <= 8'b01111100;
					mem_buffer[39:32] <= 8'b01000110;
					mem_buffer[47:40] <= 8'b01000010;
					mem_buffer[55:48] <= 8'b01000010;
					mem_buffer[63:56] <= 8'b01111100;
					end
					
			6'h0C: begin //C
					mem_buffer[7:0] <=   8'b00111110;
					mem_buffer[15:8] <=  8'b01100000;
					mem_buffer[23:16] <= 8'b01100000;
					mem_buffer[31:24] <= 8'b01100000;
					mem_buffer[39:32] <= 8'b01100000;
					mem_buffer[47:40] <= 8'b01100000;
					mem_buffer[55:48] <= 8'b01100000;
					mem_buffer[63:56] <= 8'b00111110;
					end
					
			6'h0D: begin //D
					mem_buffer[7:0] <=   8'b01111100;
					mem_buffer[15:8] <=  8'b01100010;
					mem_buffer[23:16] <= 8'b01100010;
					mem_buffer[31:24] <= 8'b01100010;
					mem_buffer[39:32] <= 8'b01100010;
					mem_buffer[47:40] <= 8'b01100010;
					mem_buffer[55:48] <= 8'b01100010;
					mem_buffer[63:56] <= 8'b01111100;
					end
					
			6'h0E: begin //E
					mem_buffer[7:0] <=   8'b00111110;
					mem_buffer[15:8] <=  8'b01100000;
					mem_buffer[23:16] <= 8'b01100000;
					mem_buffer[31:24] <= 8'b01111110;
					mem_buffer[39:32] <= 8'b01100000;
					mem_buffer[47:40] <= 8'b01100000;
					mem_buffer[55:48] <= 8'b01100000;
					mem_buffer[63:56] <= 8'b00111110;
					end
					
			6'h0F: begin //F
					mem_buffer[7:0] <=   8'b01111110;
					mem_buffer[15:8] <=  8'b01100000;
					mem_buffer[23:16] <= 8'b01100000;
					mem_buffer[31:24] <= 8'b01111110;
					mem_buffer[39:32] <= 8'b01100000;
					mem_buffer[47:40] <= 8'b01100000;
					mem_buffer[55:48] <= 8'b01100000;
					mem_buffer[63:56] <= 8'b01100000;
					end
				
			6'h10: begin //G
					mem_buffer[7:0] <=   8'b00111100;
					mem_buffer[15:8] <=  8'b01100000;
					mem_buffer[23:16] <= 8'b01100000;
					mem_buffer[31:24] <= 8'b01101110;
					mem_buffer[39:32] <= 8'b01100110;
					mem_buffer[47:40] <= 8'b01100110;
					mem_buffer[55:48] <= 8'b01100110;
					mem_buffer[63:56] <= 8'b00111100;
					end
					
			6'h11: begin //H
					mem_buffer[7:0] <=   8'b01100110;
					mem_buffer[15:8] <=  8'b01100110;
					mem_buffer[23:16] <= 8'b01100110;
					mem_buffer[31:24] <= 8'b01111110;
					mem_buffer[39:32] <= 8'b01100110;
					mem_buffer[47:40] <= 8'b01100110;
					mem_buffer[55:48] <= 8'b01100110;
					mem_buffer[63:56] <= 8'b01100110;
					end
					
			6'h12: begin //I
					mem_buffer[7:0] <=   8'b01111110;
					mem_buffer[15:8] <=  8'b00011000;
					mem_buffer[23:16] <= 8'b00011000;
					mem_buffer[31:24] <= 8'b00011000;
					mem_buffer[39:32] <= 8'b00011000;
					mem_buffer[47:40] <= 8'b00011000;
					mem_buffer[55:48] <= 8'b00011000;
					mem_buffer[63:56] <= 8'b01111110;
					end
					
			6'h13: begin //J
					mem_buffer[7:0] <=   8'b01111110;
					mem_buffer[15:8] <=  8'b00000110;
					mem_buffer[23:16] <= 8'b00000110;
					mem_buffer[31:24] <= 8'b00000110;
					mem_buffer[39:32] <= 8'b00000110;
					mem_buffer[47:40] <= 8'b00000110;
					mem_buffer[55:48] <= 8'b01100110;
					mem_buffer[63:56] <= 8'b00111100;
					end
					
			6'h14: begin //K
					mem_buffer[7:0] <=   8'b01100110;
					mem_buffer[15:8] <=  8'b01100110;
					mem_buffer[23:16] <= 8'b01101100;
					mem_buffer[31:24] <= 8'b01110000;
					mem_buffer[39:32] <= 8'b01110000;
					mem_buffer[47:40] <= 8'b01101100;
					mem_buffer[55:48] <= 8'b01100110;
					mem_buffer[63:56] <= 8'b01100110;
					end
					
			6'h15: begin //I
					mem_buffer[7:0] <=   8'b01100000;
					mem_buffer[15:8] <=  8'b01100000;
					mem_buffer[23:16] <= 8'b01100000;
					mem_buffer[31:24] <= 8'b01100000;
					mem_buffer[39:32] <= 8'b01100000;
					mem_buffer[47:40] <= 8'b01100000;
					mem_buffer[55:48] <= 8'b01100000;
					mem_buffer[63:56] <= 8'b01111110;
					end
					
			6'h16: begin //M
					mem_buffer[7:0] <=   8'b01000010;
					mem_buffer[15:8] <=  8'b01100110;
					mem_buffer[23:16] <= 8'b01011010;
					mem_buffer[31:24] <= 8'b01011010;
					mem_buffer[39:32] <= 8'b01000010;
					mem_buffer[47:40] <= 8'b01000010;
					mem_buffer[55:48] <= 8'b01000010;
					mem_buffer[63:56] <= 8'b01000010;
					end
					
			6'h17: begin //N
					mem_buffer[7:0] <=   8'b01000010;
					mem_buffer[15:8] <=  8'b01000010;
					mem_buffer[23:16] <= 8'b01100010;
					mem_buffer[31:24] <= 8'b01010010;
					mem_buffer[39:32] <= 8'b01001010;
					mem_buffer[47:40] <= 8'b01000110;
					mem_buffer[55:48] <= 8'b01000010;
					mem_buffer[63:56] <= 8'b01000010;
					end
					
			6'h18: begin //O
					mem_buffer[7:0] <=   8'b00111100;
					mem_buffer[15:8] <=  8'b01000010;
					mem_buffer[23:16] <= 8'b01000010;
					mem_buffer[31:24] <= 8'b01000010;
					mem_buffer[39:32] <= 8'b01000010;
					mem_buffer[47:40] <= 8'b01000010;
					mem_buffer[55:48] <= 8'b01000010;
					mem_buffer[63:56] <= 8'b00111100;
					end
					
			6'h19: begin //P
					mem_buffer[7:0] <=   8'b01111100;
					mem_buffer[15:8] <=  8'b01000010;
					mem_buffer[23:16] <= 8'b01000010;
					mem_buffer[31:24] <= 8'b01000010;
					mem_buffer[39:32] <= 8'b01111100;
					mem_buffer[47:40] <= 8'b01100000;
					mem_buffer[55:48] <= 8'b01100000;
					mem_buffer[63:56] <= 8'b01100000;
					end
					
			6'h1A: begin //Q
					mem_buffer[7:0] <=   8'b00111100;
					mem_buffer[15:8] <=  8'b01000010;
					mem_buffer[23:16] <= 8'b01000010;
					mem_buffer[31:24] <= 8'b01000010;
					mem_buffer[39:32] <= 8'b01000010;
					mem_buffer[47:40] <= 8'b01000010;
					mem_buffer[55:48] <= 8'b01000100;
					mem_buffer[63:56] <= 8'b00111010;
					end
					
			6'h1B: begin //R
					mem_buffer[7:0] <=   8'b00111100;
					mem_buffer[15:8] <=  8'b01000010;
					mem_buffer[23:16] <= 8'b01000010;
					mem_buffer[31:24] <= 8'b01000010;
					mem_buffer[39:32] <= 8'b01111100;
					mem_buffer[47:40] <= 8'b01011000;
					mem_buffer[55:48] <= 8'b01001100;
					mem_buffer[63:56] <= 8'b01000110;
					end
					
			6'h1C: begin //S
					mem_buffer[7:0] <=   8'b00111100;
					mem_buffer[15:8] <=  8'b01000000;
					mem_buffer[23:16] <= 8'b01000000;
					mem_buffer[31:24] <= 8'b00111100;
					mem_buffer[39:32] <= 8'b00000010;
					mem_buffer[47:40] <= 8'b00000010;
					mem_buffer[55:48] <= 8'b00000010;
					mem_buffer[63:56] <= 8'b00111100;
					end
					
			6'h1D: begin //T
					mem_buffer[7:0] <=   8'b01111110;
					mem_buffer[15:8] <=  8'b00011000;
					mem_buffer[23:16] <= 8'b00011000;
					mem_buffer[31:24] <= 8'b00011000;
					mem_buffer[39:32] <= 8'b00011000;
					mem_buffer[47:40] <= 8'b00011000;
					mem_buffer[55:48] <= 8'b00011000;
					mem_buffer[63:56] <= 8'b00011000;
					end
					
			6'h1E: begin //U
					mem_buffer[7:0] <=   8'b01000010;
					mem_buffer[15:8] <=  8'b01000010;
					mem_buffer[23:16] <= 8'b01000010;
					mem_buffer[31:24] <= 8'b01000010;
					mem_buffer[39:32] <= 8'b01000010;
					mem_buffer[47:40] <= 8'b01000010;
					mem_buffer[55:48] <= 8'b01000010;
					mem_buffer[63:56] <= 8'b00111100;
					end
					
			6'h1F: begin //V
					mem_buffer[7:0] <=   8'b01000010;
					mem_buffer[15:8] <=  8'b01000010;
					mem_buffer[23:16] <= 8'b01000010;
					mem_buffer[31:24] <= 8'b01000010;
					mem_buffer[39:32] <= 8'b01000010;
					mem_buffer[47:40] <= 8'b01000010;
					mem_buffer[55:48] <= 8'b00100100;
					mem_buffer[63:56] <= 8'b00011000;
					end
					
			6'h20: begin //W
					mem_buffer[7:0] <=   8'b01000010;
					mem_buffer[15:8] <=  8'b01000010;
					mem_buffer[23:16] <= 8'b01000010;
					mem_buffer[31:24] <= 8'b01000010;
					mem_buffer[39:32] <= 8'b01011010;
					mem_buffer[47:40] <= 8'b01011010;
					mem_buffer[55:48] <= 8'b01100110;
					mem_buffer[63:56] <= 8'b01000010;
					end
					
			6'h21: begin //X
					mem_buffer[7:0] <=   8'b01000010;
					mem_buffer[15:8] <=  8'b01000010;
					mem_buffer[23:16] <= 8'b00100100;
					mem_buffer[31:24] <= 8'b00011000;
					mem_buffer[39:32] <= 8'b00011000;
					mem_buffer[47:40] <= 8'b00100100;
					mem_buffer[55:48] <= 8'b01000010;
					mem_buffer[63:56] <= 8'b01000010;
					end
					
			6'h22: begin //Y
					mem_buffer[7:0] <=   8'b01000010;
					mem_buffer[15:8] <=  8'b01000010;
					mem_buffer[23:16] <= 8'b01000010;
					mem_buffer[31:24] <= 8'b00100100;
					mem_buffer[39:32] <= 8'b00011000;
					mem_buffer[47:40] <= 8'b00011000;
					mem_buffer[55:48] <= 8'b00011000;
					mem_buffer[63:56] <= 8'b00011000;
					end
					
			6'h23: begin //Z
					mem_buffer[7:0] <=   8'b01111110;
					mem_buffer[15:8] <=  8'b00000110;
					mem_buffer[23:16] <= 8'b00000110;
					mem_buffer[31:24] <= 8'b00001100;
					mem_buffer[39:32] <= 8'b00110000;
					mem_buffer[47:40] <= 8'b01100000;
					mem_buffer[55:48] <= 8'b01100000;
					mem_buffer[63:56] <= 8'b01111110;
					end
					
			6'h24: begin //space
					mem_buffer[7:0] <=   8'b00000000;
					mem_buffer[15:8] <=  8'b00000000;
					mem_buffer[23:16] <= 8'b00000000;
					mem_buffer[31:24] <= 8'b00000000;
					mem_buffer[39:32] <= 8'b00000000;
					mem_buffer[47:40] <= 8'b00000000;
					mem_buffer[55:48] <= 8'b00000000;
					mem_buffer[63:56] <= 8'b00000000;
					end
					
			6'h25: begin //Filled
					mem_buffer[7:0] <=   8'b11111111;
					mem_buffer[15:8] <=  8'b11111111;
					mem_buffer[23:16] <= 8'b11111111;
					mem_buffer[31:24] <= 8'b11111111;
					mem_buffer[39:32] <= 8'b11111111;
					mem_buffer[47:40] <= 8'b11111111;
					mem_buffer[55:48] <= 8'b11111111;
					mem_buffer[63:56] <= 8'b11111111;
					end
					
			6'h26: begin //-
					mem_buffer[7:0] <=   8'b00000000;
					mem_buffer[15:8] <=  8'b00000000;
					mem_buffer[23:16] <= 8'b00000000;
					mem_buffer[31:24] <= 8'b01111110;
					mem_buffer[39:32] <= 8'b00000000;
					mem_buffer[47:40] <= 8'b00000000;
					mem_buffer[55:48] <= 8'b00000000;
					mem_buffer[63:56] <= 8'b00000000;
					end
					
			6'h27: begin //:
					mem_buffer[7:0] <=   8'b00000000;
					mem_buffer[15:8] <=  8'b00011000;
					mem_buffer[23:16] <= 8'b00011000;
					mem_buffer[31:24] <= 8'b00000000;
					mem_buffer[39:32] <= 8'b00000000;
					mem_buffer[47:40] <= 8'b00011000;
					mem_buffer[55:48] <= 8'b00011000;
					mem_buffer[63:56] <= 8'b00000000;
					end
					
			6'h28: begin //.
					mem_buffer[7:0] <=   8'b00000000;
					mem_buffer[15:8] <=  8'b00000000;
					mem_buffer[23:16] <= 8'b00000000;
					mem_buffer[31:24] <= 8'b00000000;
					mem_buffer[39:32] <= 8'b00000000;
					mem_buffer[47:40] <= 8'b00000000;
					mem_buffer[55:48] <= 8'b11000000;
					mem_buffer[63:56] <= 8'b11000000;
					end
					
			default: mem_buffer <= 63'h0000000000000000;
		endcase
	endtask
endmodule	